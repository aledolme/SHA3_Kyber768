library work;
use work.keccak_globals.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity PAD_SHAKE256 is
    port(
        PADD_SHAKE256_IN : in std_logic_vector(511 downto 0);
        PADD_SHA3_OP: in std_logic_vector(1 downto 0);
        PADD_SHAKE256_OUT : out k_state
    );
end entity PAD_SHAKE256;

architecture RTL of PAD_SHAKE256 is

    signal PADD_SHAKE256_00: k_state;
    signal PADD_SHAKE256_01: k_state;

    component Keccak_2to1mux
        port(
            x      : in  k_state;
            y      : in  k_state;
            s      : in  std_logic;
            output : out k_state
        );
    end component Keccak_2to1mux;

begin

    --SHA3_OP=00
    --PADDING FOR SHAKE_256

    PADD_SHAKE256_00(0)(4)(0)<=PADD_SHAKE256_IN(56);
    PADD_SHAKE256_00(0)(4)(1)<=PADD_SHAKE256_IN(57);
    PADD_SHAKE256_00(0)(4)(2)<=PADD_SHAKE256_IN(58);
    PADD_SHAKE256_00(0)(4)(3)<=PADD_SHAKE256_IN(59);
    PADD_SHAKE256_00(0)(4)(4)<=PADD_SHAKE256_IN(60);
    PADD_SHAKE256_00(0)(4)(5)<=PADD_SHAKE256_IN(61);
    PADD_SHAKE256_00(0)(4)(6)<=PADD_SHAKE256_IN(62);
    PADD_SHAKE256_00(0)(4)(7)<=PADD_SHAKE256_IN(63);

    PADD_SHAKE256_00(0)(4)(8)<='1';
    PADD_SHAKE256_00(0)(4)(9)<='1';
    PADD_SHAKE256_00(0)(4)(10)<='1';
    PADD_SHAKE256_00(0)(4)(11)<='1';
    PADD_SHAKE256_00(0)(4)(12)<='1';
    PADD_SHAKE256_00(0)(4)(13)<='0';
    PADD_SHAKE256_00(0)(4)(14)<='0';
    PADD_SHAKE256_00(0)(4)(15)<='0';

    PADD_SHAKE256_00(0)(4)(16)<='0';
    PADD_SHAKE256_00(0)(4)(17)<='0';
    PADD_SHAKE256_00(0)(4)(18)<='0';
    PADD_SHAKE256_00(0)(4)(19)<='0';
    PADD_SHAKE256_00(0)(4)(20)<='0';
    PADD_SHAKE256_00(0)(4)(21)<='0';
    PADD_SHAKE256_00(0)(4)(22)<='0';
    PADD_SHAKE256_00(0)(4)(23)<='0';

    PADD_SHAKE256_00(0)(4)(24)<='0';
    PADD_SHAKE256_00(0)(4)(25)<='0';
    PADD_SHAKE256_00(0)(4)(26)<='0';
    PADD_SHAKE256_00(0)(4)(27)<='0';
    PADD_SHAKE256_00(0)(4)(28)<='0';
    PADD_SHAKE256_00(0)(4)(29)<='0';
    PADD_SHAKE256_00(0)(4)(30)<='0';
    PADD_SHAKE256_00(0)(4)(31)<='0';

    PADD_SHAKE256_00(0)(4)(32)<='0';
    PADD_SHAKE256_00(0)(4)(33)<='0';
    PADD_SHAKE256_00(0)(4)(34)<='0';
    PADD_SHAKE256_00(0)(4)(35)<='0';
    PADD_SHAKE256_00(0)(4)(36)<='0';
    PADD_SHAKE256_00(0)(4)(37)<='0';
    PADD_SHAKE256_00(0)(4)(38)<='0';
    PADD_SHAKE256_00(0)(4)(39)<='0';

    PADD_SHAKE256_00(0)(4)(40)<='0';
    PADD_SHAKE256_00(0)(4)(41)<='0';
    PADD_SHAKE256_00(0)(4)(42)<='0';
    PADD_SHAKE256_00(0)(4)(43)<='0';
    PADD_SHAKE256_00(0)(4)(44)<='0';
    PADD_SHAKE256_00(0)(4)(45)<='0';
    PADD_SHAKE256_00(0)(4)(46)<='0';
    PADD_SHAKE256_00(0)(4)(47)<='0';

    PADD_SHAKE256_00(0)(4)(48)<='0';
    PADD_SHAKE256_00(0)(4)(49)<='0';
    PADD_SHAKE256_00(0)(4)(50)<='0';
    PADD_SHAKE256_00(0)(4)(51)<='0';
    PADD_SHAKE256_00(0)(4)(52)<='0';
    PADD_SHAKE256_00(0)(4)(53)<='0';
    PADD_SHAKE256_00(0)(4)(54)<='0';
    PADD_SHAKE256_00(0)(4)(55)<='0';

    PADD_SHAKE256_00(0)(4)(56)<='0';
    PADD_SHAKE256_00(0)(4)(57)<='0';
    PADD_SHAKE256_00(0)(4)(58)<='0';
    PADD_SHAKE256_00(0)(4)(59)<='0';
    PADD_SHAKE256_00(0)(4)(60)<='0';
    PADD_SHAKE256_00(0)(4)(61)<='0';
    PADD_SHAKE256_00(0)(4)(62)<='0';
    PADD_SHAKE256_00(0)(4)(63)<='0';

    padd: for i in 1 to 4 generate

        PADD_SHAKE256_00(0)(4-i)(0)<=PADD_SHAKE256_IN(64+64*i-8);
        PADD_SHAKE256_00(0)(4-i)(1)<=PADD_SHAKE256_IN(64+64*i-7);
        PADD_SHAKE256_00(0)(4-i)(2)<=PADD_SHAKE256_IN(64+64*i-6);
        PADD_SHAKE256_00(0)(4-i)(3)<=PADD_SHAKE256_IN(64+64*i-5);
        PADD_SHAKE256_00(0)(4-i)(4)<=PADD_SHAKE256_IN(64+64*i-4);
        PADD_SHAKE256_00(0)(4-i)(5)<=PADD_SHAKE256_IN(64+64*i-3);
        PADD_SHAKE256_00(0)(4-i)(6)<=PADD_SHAKE256_IN(64+64*i-2);
        PADD_SHAKE256_00(0)(4-i)(7)<=PADD_SHAKE256_IN(64+64*i-1);

        PADD_SHAKE256_00(0)(4-i)(8)<=PADD_SHAKE256_IN(64+64*i-16);
        PADD_SHAKE256_00(0)(4-i)(9)<=PADD_SHAKE256_IN(64+64*i-15);
        PADD_SHAKE256_00(0)(4-i)(10)<=PADD_SHAKE256_IN(64+64*i-14);
        PADD_SHAKE256_00(0)(4-i)(11)<=PADD_SHAKE256_IN(64+64*i-13);
        PADD_SHAKE256_00(0)(4-i)(12)<=PADD_SHAKE256_IN(64+64*i-12);
        PADD_SHAKE256_00(0)(4-i)(13)<=PADD_SHAKE256_IN(64+64*i-11);
        PADD_SHAKE256_00(0)(4-i)(14)<=PADD_SHAKE256_IN(64+64*i-10);
        PADD_SHAKE256_00(0)(4-i)(15)<=PADD_SHAKE256_IN(64+64*i-9);

        PADD_SHAKE256_00(0)(4-i)(16)<=PADD_SHAKE256_IN(64+64*i-24);
        PADD_SHAKE256_00(0)(4-i)(17)<=PADD_SHAKE256_IN(64+64*i-23);
        PADD_SHAKE256_00(0)(4-i)(18)<=PADD_SHAKE256_IN(64+64*i-22);
        PADD_SHAKE256_00(0)(4-i)(19)<=PADD_SHAKE256_IN(64+64*i-21);
        PADD_SHAKE256_00(0)(4-i)(20)<=PADD_SHAKE256_IN(64+64*i-20);
        PADD_SHAKE256_00(0)(4-i)(21)<=PADD_SHAKE256_IN(64+64*i-19);
        PADD_SHAKE256_00(0)(4-i)(22)<=PADD_SHAKE256_IN(64+64*i-18);
        PADD_SHAKE256_00(0)(4-i)(23)<=PADD_SHAKE256_IN(64+64*i-17);

        PADD_SHAKE256_00(0)(4-i)(24)<=PADD_SHAKE256_IN(64+64*i-32);
        PADD_SHAKE256_00(0)(4-i)(25)<=PADD_SHAKE256_IN(64+64*i-31);
        PADD_SHAKE256_00(0)(4-i)(26)<=PADD_SHAKE256_IN(64+64*i-30);
        PADD_SHAKE256_00(0)(4-i)(27)<=PADD_SHAKE256_IN(64+64*i-29);
        PADD_SHAKE256_00(0)(4-i)(28)<=PADD_SHAKE256_IN(64+64*i-28);
        PADD_SHAKE256_00(0)(4-i)(29)<=PADD_SHAKE256_IN(64+64*i-27);
        PADD_SHAKE256_00(0)(4-i)(30)<=PADD_SHAKE256_IN(64+64*i-26);
        PADD_SHAKE256_00(0)(4-i)(31)<=PADD_SHAKE256_IN(64+64*i-25);

        PADD_SHAKE256_00(0)(4-i)(32)<=PADD_SHAKE256_IN(64+64*i-40);
        PADD_SHAKE256_00(0)(4-i)(33)<=PADD_SHAKE256_IN(64+64*i-39);
        PADD_SHAKE256_00(0)(4-i)(34)<=PADD_SHAKE256_IN(64+64*i-38);
        PADD_SHAKE256_00(0)(4-i)(35)<=PADD_SHAKE256_IN(64+64*i-37);
        PADD_SHAKE256_00(0)(4-i)(36)<=PADD_SHAKE256_IN(64+64*i-36);
        PADD_SHAKE256_00(0)(4-i)(37)<=PADD_SHAKE256_IN(64+64*i-35);
        PADD_SHAKE256_00(0)(4-i)(38)<=PADD_SHAKE256_IN(64+64*i-34);
        PADD_SHAKE256_00(0)(4-i)(39)<=PADD_SHAKE256_IN(64+64*i-33);

        PADD_SHAKE256_00(0)(4-i)(40)<=PADD_SHAKE256_IN(64+64*i-48);
        PADD_SHAKE256_00(0)(4-i)(41)<=PADD_SHAKE256_IN(64+64*i-47);
        PADD_SHAKE256_00(0)(4-i)(42)<=PADD_SHAKE256_IN(64+64*i-46);
        PADD_SHAKE256_00(0)(4-i)(43)<=PADD_SHAKE256_IN(64+64*i-45);
        PADD_SHAKE256_00(0)(4-i)(44)<=PADD_SHAKE256_IN(64+64*i-44);
        PADD_SHAKE256_00(0)(4-i)(45)<=PADD_SHAKE256_IN(64+64*i-43);
        PADD_SHAKE256_00(0)(4-i)(46)<=PADD_SHAKE256_IN(64+64*i-42);
        PADD_SHAKE256_00(0)(4-i)(47)<=PADD_SHAKE256_IN(64+64*i-41);

        PADD_SHAKE256_00(0)(4-i)(48)<=PADD_SHAKE256_IN(64+64*i-56);
        PADD_SHAKE256_00(0)(4-i)(49)<=PADD_SHAKE256_IN(64+64*i-55);
        PADD_SHAKE256_00(0)(4-i)(50)<=PADD_SHAKE256_IN(64+64*i-54);
        PADD_SHAKE256_00(0)(4-i)(51)<=PADD_SHAKE256_IN(64+64*i-53);
        PADD_SHAKE256_00(0)(4-i)(52)<=PADD_SHAKE256_IN(64+64*i-52);
        PADD_SHAKE256_00(0)(4-i)(53)<=PADD_SHAKE256_IN(64+64*i-51);
        PADD_SHAKE256_00(0)(4-i)(54)<=PADD_SHAKE256_IN(64+64*i-50);
        PADD_SHAKE256_00(0)(4-i)(55)<=PADD_SHAKE256_IN(64+64*i-49);

        PADD_SHAKE256_00(0)(4-i)(56)<=PADD_SHAKE256_IN(64+64*i-64);
        PADD_SHAKE256_00(0)(4-i)(57)<=PADD_SHAKE256_IN(64+64*i-63);
        PADD_SHAKE256_00(0)(4-i)(58)<=PADD_SHAKE256_IN(64+64*i-62);
        PADD_SHAKE256_00(0)(4-i)(59)<=PADD_SHAKE256_IN(64+64*i-61);
        PADD_SHAKE256_00(0)(4-i)(60)<=PADD_SHAKE256_IN(64+64*i-60);
        PADD_SHAKE256_00(0)(4-i)(61)<=PADD_SHAKE256_IN(64+64*i-59);
        PADD_SHAKE256_00(0)(4-i)(62)<=PADD_SHAKE256_IN(64+64*i-58);
        PADD_SHAKE256_00(0)(4-i)(63)<=PADD_SHAKE256_IN(64+64*i-57);

    end generate;


    PADD_SHAKE256_00(1)(0) <= "0000000000000000000000000000000000000000000000000000000000000000";
    PADD_SHAKE256_00(2)(0) <= "0000000000000000000000000000000000000000000000000000000000000000";
    PADD_SHAKE256_00(3)(0) <= "0000000000000000000000000000000000000000000000000000000000000000";
    PADD_SHAKE256_00(4)(0) <= "0000000000000000000000000000000000000000000000000000000000000000";

    PADD_SHAKE256_00(1)(1) <= "0000000000000000000000000000000000000000000000000000000000000000";
    PADD_SHAKE256_00(2)(1) <= "0000000000000000000000000000000000000000000000000000000000000000";
    PADD_SHAKE256_00(3)(1) <= "1000000000000000000000000000000000000000000000000000000000000000";
    PADD_SHAKE256_00(4)(1) <= "0000000000000000000000000000000000000000000000000000000000000000";

    PADD_SHAKE256_00(1)(2) <= "0000000000000000000000000000000000000000000000000000000000000000";
    PADD_SHAKE256_00(2)(2) <= "0000000000000000000000000000000000000000000000000000000000000000";
    PADD_SHAKE256_00(3)(2) <= "0000000000000000000000000000000000000000000000000000000000000000";
    PADD_SHAKE256_00(4)(2) <= "0000000000000000000000000000000000000000000000000000000000000000";

    PADD_SHAKE256_00(1)(3) <= "0000000000000000000000000000000000000000000000000000000000000000";
    PADD_SHAKE256_00(2)(3) <= "0000000000000000000000000000000000000000000000000000000000000000";
    PADD_SHAKE256_00(3)(3) <= "0000000000000000000000000000000000000000000000000000000000000000";
    PADD_SHAKE256_00(4)(3) <= "0000000000000000000000000000000000000000000000000000000000000000";

    PADD_SHAKE256_00(1)(4) <= "0000000000000000000000000000000000000000000000000000000000000000";
    PADD_SHAKE256_00(2)(4) <= "0000000000000000000000000000000000000000000000000000000000000000";
    PADD_SHAKE256_00(3)(4) <= "0000000000000000000000000000000000000000000000000000000000000000";
    PADD_SHAKE256_00(4)(4) <= "0000000000000000000000000000000000000000000000000000000000000000";



    --SHAE_OP=01
    --PADDING FOR SHAKE_256

    padd01: for i in 1 to 5 generate

        PADD_SHAKE256_01(0)(5-i)(0)<=PADD_SHAKE256_IN(192+64*i-8);
        PADD_SHAKE256_01(0)(5-i)(1)<=PADD_SHAKE256_IN(192+64*i-7);
        PADD_SHAKE256_01(0)(5-i)(2)<=PADD_SHAKE256_IN(192+64*i-6);
        PADD_SHAKE256_01(0)(5-i)(3)<=PADD_SHAKE256_IN(192+64*i-5);
        PADD_SHAKE256_01(0)(5-i)(4)<=PADD_SHAKE256_IN(192+64*i-4);
        PADD_SHAKE256_01(0)(5-i)(5)<=PADD_SHAKE256_IN(192+64*i-3);
        PADD_SHAKE256_01(0)(5-i)(6)<=PADD_SHAKE256_IN(192+64*i-2);
        PADD_SHAKE256_01(0)(5-i)(7)<=PADD_SHAKE256_IN(192+64*i-1);

        PADD_SHAKE256_01(0)(5-i)(8)<=PADD_SHAKE256_IN(192+64*i-16);
        PADD_SHAKE256_01(0)(5-i)(9)<=PADD_SHAKE256_IN(192+64*i-15);
        PADD_SHAKE256_01(0)(5-i)(10)<=PADD_SHAKE256_IN(192+64*i-14);
        PADD_SHAKE256_01(0)(5-i)(11)<=PADD_SHAKE256_IN(192+64*i-13);
        PADD_SHAKE256_01(0)(5-i)(12)<=PADD_SHAKE256_IN(192+64*i-12);
        PADD_SHAKE256_01(0)(5-i)(13)<=PADD_SHAKE256_IN(192+64*i-11);
        PADD_SHAKE256_01(0)(5-i)(14)<=PADD_SHAKE256_IN(192+64*i-10);
        PADD_SHAKE256_01(0)(5-i)(15)<=PADD_SHAKE256_IN(192+64*i-9);

        PADD_SHAKE256_01(0)(5-i)(16)<=PADD_SHAKE256_IN(192+64*i-24);
        PADD_SHAKE256_01(0)(5-i)(17)<=PADD_SHAKE256_IN(192+64*i-23);
        PADD_SHAKE256_01(0)(5-i)(18)<=PADD_SHAKE256_IN(192+64*i-22);
        PADD_SHAKE256_01(0)(5-i)(19)<=PADD_SHAKE256_IN(192+64*i-21);
        PADD_SHAKE256_01(0)(5-i)(20)<=PADD_SHAKE256_IN(192+64*i-20);
        PADD_SHAKE256_01(0)(5-i)(21)<=PADD_SHAKE256_IN(192+64*i-19);
        PADD_SHAKE256_01(0)(5-i)(22)<=PADD_SHAKE256_IN(192+64*i-18);
        PADD_SHAKE256_01(0)(5-i)(23)<=PADD_SHAKE256_IN(192+64*i-17);

        PADD_SHAKE256_01(0)(5-i)(24)<=PADD_SHAKE256_IN(192+64*i-32);
        PADD_SHAKE256_01(0)(5-i)(25)<=PADD_SHAKE256_IN(192+64*i-31);
        PADD_SHAKE256_01(0)(5-i)(26)<=PADD_SHAKE256_IN(192+64*i-30);
        PADD_SHAKE256_01(0)(5-i)(27)<=PADD_SHAKE256_IN(192+64*i-29);
        PADD_SHAKE256_01(0)(5-i)(28)<=PADD_SHAKE256_IN(192+64*i-28);
        PADD_SHAKE256_01(0)(5-i)(29)<=PADD_SHAKE256_IN(192+64*i-27);
        PADD_SHAKE256_01(0)(5-i)(30)<=PADD_SHAKE256_IN(192+64*i-26);
        PADD_SHAKE256_01(0)(5-i)(31)<=PADD_SHAKE256_IN(192+64*i-25);

        PADD_SHAKE256_01(0)(5-i)(32)<=PADD_SHAKE256_IN(192+64*i-40);
        PADD_SHAKE256_01(0)(5-i)(33)<=PADD_SHAKE256_IN(192+64*i-39);
        PADD_SHAKE256_01(0)(5-i)(34)<=PADD_SHAKE256_IN(192+64*i-38);
        PADD_SHAKE256_01(0)(5-i)(35)<=PADD_SHAKE256_IN(192+64*i-37);
        PADD_SHAKE256_01(0)(5-i)(36)<=PADD_SHAKE256_IN(192+64*i-36);
        PADD_SHAKE256_01(0)(5-i)(37)<=PADD_SHAKE256_IN(192+64*i-35);
        PADD_SHAKE256_01(0)(5-i)(38)<=PADD_SHAKE256_IN(192+64*i-34);
        PADD_SHAKE256_01(0)(5-i)(39)<=PADD_SHAKE256_IN(192+64*i-33);

        PADD_SHAKE256_01(0)(5-i)(40)<=PADD_SHAKE256_IN(192+64*i-48);
        PADD_SHAKE256_01(0)(5-i)(41)<=PADD_SHAKE256_IN(192+64*i-47);
        PADD_SHAKE256_01(0)(5-i)(42)<=PADD_SHAKE256_IN(192+64*i-46);
        PADD_SHAKE256_01(0)(5-i)(43)<=PADD_SHAKE256_IN(192+64*i-45);
        PADD_SHAKE256_01(0)(5-i)(44)<=PADD_SHAKE256_IN(192+64*i-44);
        PADD_SHAKE256_01(0)(5-i)(45)<=PADD_SHAKE256_IN(192+64*i-43);
        PADD_SHAKE256_01(0)(5-i)(46)<=PADD_SHAKE256_IN(192+64*i-42);
        PADD_SHAKE256_01(0)(5-i)(47)<=PADD_SHAKE256_IN(192+64*i-41);

        PADD_SHAKE256_01(0)(5-i)(48)<=PADD_SHAKE256_IN(192+64*i-56);
        PADD_SHAKE256_01(0)(5-i)(49)<=PADD_SHAKE256_IN(192+64*i-55);
        PADD_SHAKE256_01(0)(5-i)(50)<=PADD_SHAKE256_IN(192+64*i-54);
        PADD_SHAKE256_01(0)(5-i)(51)<=PADD_SHAKE256_IN(192+64*i-53);
        PADD_SHAKE256_01(0)(5-i)(52)<=PADD_SHAKE256_IN(192+64*i-52);
        PADD_SHAKE256_01(0)(5-i)(53)<=PADD_SHAKE256_IN(192+64*i-51);
        PADD_SHAKE256_01(0)(5-i)(54)<=PADD_SHAKE256_IN(192+64*i-50);
        PADD_SHAKE256_01(0)(5-i)(55)<=PADD_SHAKE256_IN(192+64*i-49);

        PADD_SHAKE256_01(0)(5-i)(56)<=PADD_SHAKE256_IN(192+64*i-64);
        PADD_SHAKE256_01(0)(5-i)(57)<=PADD_SHAKE256_IN(192+64*i-63);
        PADD_SHAKE256_01(0)(5-i)(58)<=PADD_SHAKE256_IN(192+64*i-62);
        PADD_SHAKE256_01(0)(5-i)(59)<=PADD_SHAKE256_IN(192+64*i-61);
        PADD_SHAKE256_01(0)(5-i)(60)<=PADD_SHAKE256_IN(192+64*i-60);
        PADD_SHAKE256_01(0)(5-i)(61)<=PADD_SHAKE256_IN(192+64*i-59);
        PADD_SHAKE256_01(0)(5-i)(62)<=PADD_SHAKE256_IN(192+64*i-58);
        PADD_SHAKE256_01(0)(5-i)(63)<=PADD_SHAKE256_IN(192+64*i-57);

    end generate;

    padd03: for i in 1 to 3 generate

        PADD_SHAKE256_01(1)(3-i)(0)<=PADD_SHAKE256_IN(64*i-8);
        PADD_SHAKE256_01(1)(3-i)(1)<=PADD_SHAKE256_IN(64*i-7);
        PADD_SHAKE256_01(1)(3-i)(2)<=PADD_SHAKE256_IN(64*i-6);
        PADD_SHAKE256_01(1)(3-i)(3)<=PADD_SHAKE256_IN(64*i-5);
        PADD_SHAKE256_01(1)(3-i)(4)<=PADD_SHAKE256_IN(64*i-4);
        PADD_SHAKE256_01(1)(3-i)(5)<=PADD_SHAKE256_IN(64*i-3);
        PADD_SHAKE256_01(1)(3-i)(6)<=PADD_SHAKE256_IN(64*i-2);
        PADD_SHAKE256_01(1)(3-i)(7)<=PADD_SHAKE256_IN(64*i-1);

        PADD_SHAKE256_01(1)(3-i)(8)<=PADD_SHAKE256_IN(64*i-16);
        PADD_SHAKE256_01(1)(3-i)(9)<=PADD_SHAKE256_IN(64*i-15);
        PADD_SHAKE256_01(1)(3-i)(10)<=PADD_SHAKE256_IN(64*i-14);
        PADD_SHAKE256_01(1)(3-i)(11)<=PADD_SHAKE256_IN(64*i-13);
        PADD_SHAKE256_01(1)(3-i)(12)<=PADD_SHAKE256_IN(64*i-12);
        PADD_SHAKE256_01(1)(3-i)(13)<=PADD_SHAKE256_IN(64*i-11);
        PADD_SHAKE256_01(1)(3-i)(14)<=PADD_SHAKE256_IN(64*i-10);
        PADD_SHAKE256_01(1)(3-i)(15)<=PADD_SHAKE256_IN(64*i-9);

        PADD_SHAKE256_01(1)(3-i)(16)<=PADD_SHAKE256_IN(64*i-24);
        PADD_SHAKE256_01(1)(3-i)(17)<=PADD_SHAKE256_IN(64*i-23);
        PADD_SHAKE256_01(1)(3-i)(18)<=PADD_SHAKE256_IN(64*i-22);
        PADD_SHAKE256_01(1)(3-i)(19)<=PADD_SHAKE256_IN(64*i-21);
        PADD_SHAKE256_01(1)(3-i)(20)<=PADD_SHAKE256_IN(64*i-20);
        PADD_SHAKE256_01(1)(3-i)(21)<=PADD_SHAKE256_IN(64*i-19);
        PADD_SHAKE256_01(1)(3-i)(22)<=PADD_SHAKE256_IN(64*i-18);
        PADD_SHAKE256_01(1)(3-i)(23)<=PADD_SHAKE256_IN(64*i-17);

        PADD_SHAKE256_01(1)(3-i)(24)<=PADD_SHAKE256_IN(64*i-32);
        PADD_SHAKE256_01(1)(3-i)(25)<=PADD_SHAKE256_IN(64*i-31);
        PADD_SHAKE256_01(1)(3-i)(26)<=PADD_SHAKE256_IN(64*i-30);
        PADD_SHAKE256_01(1)(3-i)(27)<=PADD_SHAKE256_IN(64*i-29);
        PADD_SHAKE256_01(1)(3-i)(28)<=PADD_SHAKE256_IN(64*i-28);
        PADD_SHAKE256_01(1)(3-i)(29)<=PADD_SHAKE256_IN(64*i-27);
        PADD_SHAKE256_01(1)(3-i)(30)<=PADD_SHAKE256_IN(64*i-26);
        PADD_SHAKE256_01(1)(3-i)(31)<=PADD_SHAKE256_IN(64*i-25);

        PADD_SHAKE256_01(1)(3-i)(32)<=PADD_SHAKE256_IN(64*i-40);
        PADD_SHAKE256_01(1)(3-i)(33)<=PADD_SHAKE256_IN(64*i-39);
        PADD_SHAKE256_01(1)(3-i)(34)<=PADD_SHAKE256_IN(64*i-38);
        PADD_SHAKE256_01(1)(3-i)(35)<=PADD_SHAKE256_IN(64*i-37);
        PADD_SHAKE256_01(1)(3-i)(36)<=PADD_SHAKE256_IN(64*i-36);
        PADD_SHAKE256_01(1)(3-i)(37)<=PADD_SHAKE256_IN(64*i-35);
        PADD_SHAKE256_01(1)(3-i)(38)<=PADD_SHAKE256_IN(64*i-34);
        PADD_SHAKE256_01(1)(3-i)(39)<=PADD_SHAKE256_IN(64*i-33);

        PADD_SHAKE256_01(1)(3-i)(40)<=PADD_SHAKE256_IN(64*i-48);
        PADD_SHAKE256_01(1)(3-i)(41)<=PADD_SHAKE256_IN(64*i-47);
        PADD_SHAKE256_01(1)(3-i)(42)<=PADD_SHAKE256_IN(64*i-46);
        PADD_SHAKE256_01(1)(3-i)(43)<=PADD_SHAKE256_IN(64*i-45);
        PADD_SHAKE256_01(1)(3-i)(44)<=PADD_SHAKE256_IN(64*i-44);
        PADD_SHAKE256_01(1)(3-i)(45)<=PADD_SHAKE256_IN(64*i-43);
        PADD_SHAKE256_01(1)(3-i)(46)<=PADD_SHAKE256_IN(64*i-42);
        PADD_SHAKE256_01(1)(3-i)(47)<=PADD_SHAKE256_IN(64*i-41);

        PADD_SHAKE256_01(1)(3-i)(48)<=PADD_SHAKE256_IN(64*i-56);
        PADD_SHAKE256_01(1)(3-i)(49)<=PADD_SHAKE256_IN(64*i-55);
        PADD_SHAKE256_01(1)(3-i)(50)<=PADD_SHAKE256_IN(64*i-54);
        PADD_SHAKE256_01(1)(3-i)(51)<=PADD_SHAKE256_IN(64*i-53);
        PADD_SHAKE256_01(1)(3-i)(52)<=PADD_SHAKE256_IN(64*i-52);
        PADD_SHAKE256_01(1)(3-i)(53)<=PADD_SHAKE256_IN(64*i-51);
        PADD_SHAKE256_01(1)(3-i)(54)<=PADD_SHAKE256_IN(64*i-50);
        PADD_SHAKE256_01(1)(3-i)(55)<=PADD_SHAKE256_IN(64*i-49);

        PADD_SHAKE256_01(1)(3-i)(56)<=PADD_SHAKE256_IN(64*i-64);
        PADD_SHAKE256_01(1)(3-i)(57)<=PADD_SHAKE256_IN(64*i-63);
        PADD_SHAKE256_01(1)(3-i)(58)<=PADD_SHAKE256_IN(64*i-62);
        PADD_SHAKE256_01(1)(3-i)(59)<=PADD_SHAKE256_IN(64*i-61);
        PADD_SHAKE256_01(1)(3-i)(60)<=PADD_SHAKE256_IN(64*i-60);
        PADD_SHAKE256_01(1)(3-i)(61)<=PADD_SHAKE256_IN(64*i-59);
        PADD_SHAKE256_01(1)(3-i)(62)<=PADD_SHAKE256_IN(64*i-58);
        PADD_SHAKE256_01(1)(3-i)(63)<=PADD_SHAKE256_IN(64*i-57);

    end generate;

    PADD_SHAKE256_01(2)(0) <= "0000000000000000000000000000000000000000000000000000000000000000";
    PADD_SHAKE256_01(3)(0) <= "0000000000000000000000000000000000000000000000000000000000000000";
    PADD_SHAKE256_01(4)(0) <= "0000000000000000000000000000000000000000000000000000000000000000";

    PADD_SHAKE256_01(2)(1) <= "0000000000000000000000000000000000000000000000000000000000000000";
    PADD_SHAKE256_01(3)(1) <= "1000000000000000000000000000000000000000000000000000000000000000";
    PADD_SHAKE256_01(4)(1) <= "0000000000000000000000000000000000000000000000000000000000000000";

    PADD_SHAKE256_01(2)(2) <= "0000000000000000000000000000000000000000000000000000000000000000";
    PADD_SHAKE256_01(3)(2) <= "0000000000000000000000000000000000000000000000000000000000000000";
    PADD_SHAKE256_01(4)(2) <= "0000000000000000000000000000000000000000000000000000000000000000";

    PADD_SHAKE256_01(1)(3) <= "0000000000000000000000000000000000000000000000000000000000011111";
    PADD_SHAKE256_01(2)(3) <= "0000000000000000000000000000000000000000000000000000000000000000";
    PADD_SHAKE256_01(3)(3) <= "0000000000000000000000000000000000000000000000000000000000000000";
    PADD_SHAKE256_01(4)(3) <= "0000000000000000000000000000000000000000000000000000000000000000";

    PADD_SHAKE256_01(1)(4) <= "0000000000000000000000000000000000000000000000000000000000000000";
    PADD_SHAKE256_01(2)(4) <= "0000000000000000000000000000000000000000000000000000000000000000";
    PADD_SHAKE256_01(3)(4) <= "0000000000000000000000000000000000000000000000000000000000000000";
    PADD_SHAKE256_01(4)(4) <= "0000000000000000000000000000000000000000000000000000000000000000";


    i_mux_SHAKE256: Keccak_2to1mux
        port map(
            x      => PADD_SHAKE256_00,
            y      => PADD_SHAKE256_01,
            s      => PADD_SHA3_OP(0),
            output => PADD_SHAKE256_OUT
        );

end architecture RTL;
