library work;
use work.keccak_globals.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity PAD_SHAKE128 is
    port(
        PADD_SHAKE128_IN : in std_logic_vector(271 downto 0);
        PADD_SHAKE128_OUT : out k_state
    );
end entity PAD_SHAKE128;

architecture RTL of PAD_SHAKE128 is

begin

    --SHAE_OP=00
    --PADDING FOR SHAKE_128

    PADD_SHAKE128_OUT(0)(4)(0)<=PADD_SHAKE128_IN(8);
    PADD_SHAKE128_OUT(0)(4)(1)<=PADD_SHAKE128_IN(9);
    PADD_SHAKE128_OUT(0)(4)(2)<=PADD_SHAKE128_IN(10);
    PADD_SHAKE128_OUT(0)(4)(3)<=PADD_SHAKE128_IN(11);
    PADD_SHAKE128_OUT(0)(4)(4)<=PADD_SHAKE128_IN(12);
    PADD_SHAKE128_OUT(0)(4)(5)<=PADD_SHAKE128_IN(13);
    PADD_SHAKE128_OUT(0)(4)(6)<=PADD_SHAKE128_IN(14);
    PADD_SHAKE128_OUT(0)(4)(7)<=PADD_SHAKE128_IN(15);

    PADD_SHAKE128_OUT(0)(4)(8)<=PADD_SHAKE128_IN(0);
    PADD_SHAKE128_OUT(0)(4)(9)<=PADD_SHAKE128_IN(1);
    PADD_SHAKE128_OUT(0)(4)(10)<=PADD_SHAKE128_IN(2);
    PADD_SHAKE128_OUT(0)(4)(11)<=PADD_SHAKE128_IN(3);
    PADD_SHAKE128_OUT(0)(4)(12)<=PADD_SHAKE128_IN(4);
    PADD_SHAKE128_OUT(0)(4)(13)<=PADD_SHAKE128_IN(5);
    PADD_SHAKE128_OUT(0)(4)(14)<=PADD_SHAKE128_IN(6);
    PADD_SHAKE128_OUT(0)(4)(15)<=PADD_SHAKE128_IN(7);

    PADD_SHAKE128_OUT(0)(4)(16)<='1';
    PADD_SHAKE128_OUT(0)(4)(17)<='1';
    PADD_SHAKE128_OUT(0)(4)(18)<='1';
    PADD_SHAKE128_OUT(0)(4)(19)<='1';
    PADD_SHAKE128_OUT(0)(4)(20)<='1';
    PADD_SHAKE128_OUT(0)(4)(21)<='0';
    PADD_SHAKE128_OUT(0)(4)(22)<='0';
    PADD_SHAKE128_OUT(0)(4)(23)<='0';

    PADD_SHAKE128_OUT(0)(4)(24)<='0';
    PADD_SHAKE128_OUT(0)(4)(25)<='0';
    PADD_SHAKE128_OUT(0)(4)(26)<='0';
    PADD_SHAKE128_OUT(0)(4)(27)<='0';
    PADD_SHAKE128_OUT(0)(4)(28)<='0';
    PADD_SHAKE128_OUT(0)(4)(29)<='0';
    PADD_SHAKE128_OUT(0)(4)(30)<='0';
    PADD_SHAKE128_OUT(0)(4)(31)<='0';

    PADD_SHAKE128_OUT(0)(4)(32)<='0';
    PADD_SHAKE128_OUT(0)(4)(33)<='0';
    PADD_SHAKE128_OUT(0)(4)(34)<='0';
    PADD_SHAKE128_OUT(0)(4)(35)<='0';
    PADD_SHAKE128_OUT(0)(4)(36)<='0';
    PADD_SHAKE128_OUT(0)(4)(37)<='0';
    PADD_SHAKE128_OUT(0)(4)(38)<='0';
    PADD_SHAKE128_OUT(0)(4)(39)<='0';

    PADD_SHAKE128_OUT(0)(4)(40)<='0';
    PADD_SHAKE128_OUT(0)(4)(41)<='0';
    PADD_SHAKE128_OUT(0)(4)(42)<='0';
    PADD_SHAKE128_OUT(0)(4)(43)<='0';
    PADD_SHAKE128_OUT(0)(4)(44)<='0';
    PADD_SHAKE128_OUT(0)(4)(45)<='0';
    PADD_SHAKE128_OUT(0)(4)(46)<='0';
    PADD_SHAKE128_OUT(0)(4)(47)<='0';

    PADD_SHAKE128_OUT(0)(4)(48)<='0';
    PADD_SHAKE128_OUT(0)(4)(49)<='0';
    PADD_SHAKE128_OUT(0)(4)(50)<='0';
    PADD_SHAKE128_OUT(0)(4)(51)<='0';
    PADD_SHAKE128_OUT(0)(4)(52)<='0';
    PADD_SHAKE128_OUT(0)(4)(53)<='0';
    PADD_SHAKE128_OUT(0)(4)(54)<='0';
    PADD_SHAKE128_OUT(0)(4)(55)<='0';

    PADD_SHAKE128_OUT(0)(4)(56)<='0';
    PADD_SHAKE128_OUT(0)(4)(57)<='0';
    PADD_SHAKE128_OUT(0)(4)(58)<='0';
    PADD_SHAKE128_OUT(0)(4)(59)<='0';
    PADD_SHAKE128_OUT(0)(4)(60)<='0';
    PADD_SHAKE128_OUT(0)(4)(61)<='0';
    PADD_SHAKE128_OUT(0)(4)(62)<='0';
    PADD_SHAKE128_OUT(0)(4)(63)<='0';

    padd: for i in 1 to 4 generate

        PADD_SHAKE128_OUT(0)(4-i)(0)<=PADD_SHAKE128_IN(16+64*i-8);
        PADD_SHAKE128_OUT(0)(4-i)(1)<=PADD_SHAKE128_IN(16+64*i-7);
        PADD_SHAKE128_OUT(0)(4-i)(2)<=PADD_SHAKE128_IN(16+64*i-6);
        PADD_SHAKE128_OUT(0)(4-i)(3)<=PADD_SHAKE128_IN(16+64*i-5);
        PADD_SHAKE128_OUT(0)(4-i)(4)<=PADD_SHAKE128_IN(16+64*i-4);
        PADD_SHAKE128_OUT(0)(4-i)(5)<=PADD_SHAKE128_IN(16+64*i-3);
        PADD_SHAKE128_OUT(0)(4-i)(6)<=PADD_SHAKE128_IN(16+64*i-2);
        PADD_SHAKE128_OUT(0)(4-i)(7)<=PADD_SHAKE128_IN(16+64*i-1);

        PADD_SHAKE128_OUT(0)(4-i)(8)<=PADD_SHAKE128_IN(16+64*i-16);
        PADD_SHAKE128_OUT(0)(4-i)(9)<=PADD_SHAKE128_IN(16+64*i-15);
        PADD_SHAKE128_OUT(0)(4-i)(10)<=PADD_SHAKE128_IN(16+64*i-14);
        PADD_SHAKE128_OUT(0)(4-i)(11)<=PADD_SHAKE128_IN(16+64*i-13);
        PADD_SHAKE128_OUT(0)(4-i)(12)<=PADD_SHAKE128_IN(16+64*i-12);
        PADD_SHAKE128_OUT(0)(4-i)(13)<=PADD_SHAKE128_IN(16+64*i-11);
        PADD_SHAKE128_OUT(0)(4-i)(14)<=PADD_SHAKE128_IN(16+64*i-10);
        PADD_SHAKE128_OUT(0)(4-i)(15)<=PADD_SHAKE128_IN(16+64*i-9);

        PADD_SHAKE128_OUT(0)(4-i)(16)<=PADD_SHAKE128_IN(16+64*i-24);
        PADD_SHAKE128_OUT(0)(4-i)(17)<=PADD_SHAKE128_IN(16+64*i-23);
        PADD_SHAKE128_OUT(0)(4-i)(18)<=PADD_SHAKE128_IN(16+64*i-22);
        PADD_SHAKE128_OUT(0)(4-i)(19)<=PADD_SHAKE128_IN(16+64*i-21);
        PADD_SHAKE128_OUT(0)(4-i)(20)<=PADD_SHAKE128_IN(16+64*i-20);
        PADD_SHAKE128_OUT(0)(4-i)(21)<=PADD_SHAKE128_IN(16+64*i-19);
        PADD_SHAKE128_OUT(0)(4-i)(22)<=PADD_SHAKE128_IN(16+64*i-18);
        PADD_SHAKE128_OUT(0)(4-i)(23)<=PADD_SHAKE128_IN(16+64*i-17);

        PADD_SHAKE128_OUT(0)(4-i)(24)<=PADD_SHAKE128_IN(16+64*i-32);
        PADD_SHAKE128_OUT(0)(4-i)(25)<=PADD_SHAKE128_IN(16+64*i-31);
        PADD_SHAKE128_OUT(0)(4-i)(26)<=PADD_SHAKE128_IN(16+64*i-30);
        PADD_SHAKE128_OUT(0)(4-i)(27)<=PADD_SHAKE128_IN(16+64*i-29);
        PADD_SHAKE128_OUT(0)(4-i)(28)<=PADD_SHAKE128_IN(16+64*i-28);
        PADD_SHAKE128_OUT(0)(4-i)(29)<=PADD_SHAKE128_IN(16+64*i-27);
        PADD_SHAKE128_OUT(0)(4-i)(30)<=PADD_SHAKE128_IN(16+64*i-26);
        PADD_SHAKE128_OUT(0)(4-i)(31)<=PADD_SHAKE128_IN(16+64*i-25);

        PADD_SHAKE128_OUT(0)(4-i)(32)<=PADD_SHAKE128_IN(16+64*i-40);
        PADD_SHAKE128_OUT(0)(4-i)(33)<=PADD_SHAKE128_IN(16+64*i-39);
        PADD_SHAKE128_OUT(0)(4-i)(34)<=PADD_SHAKE128_IN(16+64*i-38);
        PADD_SHAKE128_OUT(0)(4-i)(35)<=PADD_SHAKE128_IN(16+64*i-37);
        PADD_SHAKE128_OUT(0)(4-i)(36)<=PADD_SHAKE128_IN(16+64*i-36);
        PADD_SHAKE128_OUT(0)(4-i)(37)<=PADD_SHAKE128_IN(16+64*i-35);
        PADD_SHAKE128_OUT(0)(4-i)(38)<=PADD_SHAKE128_IN(16+64*i-34);
        PADD_SHAKE128_OUT(0)(4-i)(39)<=PADD_SHAKE128_IN(16+64*i-33);

        PADD_SHAKE128_OUT(0)(4-i)(40)<=PADD_SHAKE128_IN(16+64*i-48);
        PADD_SHAKE128_OUT(0)(4-i)(41)<=PADD_SHAKE128_IN(16+64*i-47);
        PADD_SHAKE128_OUT(0)(4-i)(42)<=PADD_SHAKE128_IN(16+64*i-46);
        PADD_SHAKE128_OUT(0)(4-i)(43)<=PADD_SHAKE128_IN(16+64*i-45);
        PADD_SHAKE128_OUT(0)(4-i)(44)<=PADD_SHAKE128_IN(16+64*i-44);
        PADD_SHAKE128_OUT(0)(4-i)(45)<=PADD_SHAKE128_IN(16+64*i-43);
        PADD_SHAKE128_OUT(0)(4-i)(46)<=PADD_SHAKE128_IN(16+64*i-42);
        PADD_SHAKE128_OUT(0)(4-i)(47)<=PADD_SHAKE128_IN(16+64*i-41);

        PADD_SHAKE128_OUT(0)(4-i)(48)<=PADD_SHAKE128_IN(16+64*i-56);
        PADD_SHAKE128_OUT(0)(4-i)(49)<=PADD_SHAKE128_IN(16+64*i-55);
        PADD_SHAKE128_OUT(0)(4-i)(50)<=PADD_SHAKE128_IN(16+64*i-54);
        PADD_SHAKE128_OUT(0)(4-i)(51)<=PADD_SHAKE128_IN(16+64*i-53);
        PADD_SHAKE128_OUT(0)(4-i)(52)<=PADD_SHAKE128_IN(16+64*i-52);
        PADD_SHAKE128_OUT(0)(4-i)(53)<=PADD_SHAKE128_IN(16+64*i-51);
        PADD_SHAKE128_OUT(0)(4-i)(54)<=PADD_SHAKE128_IN(16+64*i-50);
        PADD_SHAKE128_OUT(0)(4-i)(55)<=PADD_SHAKE128_IN(16+64*i-49);

        PADD_SHAKE128_OUT(0)(4-i)(56)<=PADD_SHAKE128_IN(16+64*i-64);
        PADD_SHAKE128_OUT(0)(4-i)(57)<=PADD_SHAKE128_IN(16+64*i-63);
        PADD_SHAKE128_OUT(0)(4-i)(58)<=PADD_SHAKE128_IN(16+64*i-62);
        PADD_SHAKE128_OUT(0)(4-i)(59)<=PADD_SHAKE128_IN(16+64*i-61);
        PADD_SHAKE128_OUT(0)(4-i)(60)<=PADD_SHAKE128_IN(16+64*i-60);
        PADD_SHAKE128_OUT(0)(4-i)(61)<=PADD_SHAKE128_IN(16+64*i-59);
        PADD_SHAKE128_OUT(0)(4-i)(62)<=PADD_SHAKE128_IN(16+64*i-58);
        PADD_SHAKE128_OUT(0)(4-i)(63)<=PADD_SHAKE128_IN(16+64*i-57);

    end generate;



    PADD_SHAKE128_OUT(1)(0) <= "0000000000000000000000000000000000000000000000000000000000000000";
    PADD_SHAKE128_OUT(2)(0) <= "0000000000000000000000000000000000000000000000000000000000000000";
    PADD_SHAKE128_OUT(3)(0) <= "0000000000000000000000000000000000000000000000000000000000000000";
    PADD_SHAKE128_OUT(4)(0) <= "1000000000000000000000000000000000000000000000000000000000000000";

    PADD_SHAKE128_OUT(1)(1) <= "0000000000000000000000000000000000000000000000000000000000000000";
    PADD_SHAKE128_OUT(2)(1) <= "0000000000000000000000000000000000000000000000000000000000000000";
    PADD_SHAKE128_OUT(3)(1) <= "0000000000000000000000000000000000000000000000000000000000000000";
    PADD_SHAKE128_OUT(4)(1) <= "0000000000000000000000000000000000000000000000000000000000000000";

    PADD_SHAKE128_OUT(1)(2) <= "0000000000000000000000000000000000000000000000000000000000000000";
    PADD_SHAKE128_OUT(2)(2) <= "0000000000000000000000000000000000000000000000000000000000000000";
    PADD_SHAKE128_OUT(3)(2) <= "0000000000000000000000000000000000000000000000000000000000000000";
    PADD_SHAKE128_OUT(4)(2) <= "0000000000000000000000000000000000000000000000000000000000000000";

    PADD_SHAKE128_OUT(1)(3) <= "0000000000000000000000000000000000000000000000000000000000000000";
    PADD_SHAKE128_OUT(2)(3) <= "0000000000000000000000000000000000000000000000000000000000000000";
    PADD_SHAKE128_OUT(3)(3) <= "0000000000000000000000000000000000000000000000000000000000000000";
    PADD_SHAKE128_OUT(4)(3) <= "0000000000000000000000000000000000000000000000000000000000000000";

    PADD_SHAKE128_OUT(1)(4) <= "0000000000000000000000000000000000000000000000000000000000000000";
    PADD_SHAKE128_OUT(2)(4) <= "0000000000000000000000000000000000000000000000000000000000000000";
    PADD_SHAKE128_OUT(3)(4) <= "0000000000000000000000000000000000000000000000000000000000000000";
    PADD_SHAKE128_OUT(4)(4) <= "0000000000000000000000000000000000000000000000000000000000000000";




end architecture RTL;
